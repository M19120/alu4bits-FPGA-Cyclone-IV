library verilog;
use verilog.vl_types.all;
entity alu_4bits_vlg_vec_tst is
end alu_4bits_vlg_vec_tst;
